package definitions is
constant N : integer := 6;
constant M : integer := 3;
constant W_CONTROL : integer := 9;
constant W_STATUS : integer := 2;
-- Control Constants
-- <DEFINE>
-- constant W_CONTROL : integer := <DEFINE>; -- Control vector width
-- Status Constants
-- <DEFINE>
-- constant W_STATUS : integer := <DEFINE>; -- Status vector width
end package definitions;